`include"./qmult.sv"
module tb();
logic [255:0] n1,n2;
logic [255:0]r;
logic f;
qmult m(1'b1,n1,n1,r,f);

initial begin
    $monitor("%h.%h^2 =  %h.%h\n",n1[255:16],n1[15:0],r[255:16],r[15:0]);
    #1 n1 = 256'b0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000001_1110000000000000;
    #1 n1 = r;
    #1 n1 = r;
    #1 n1 = r;
    #1 n1 = r;
    #1 n1 = r;
    #1 n1 = r;

end
endmodule
//00000000000000000